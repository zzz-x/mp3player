module Char_Set(
	 input[4:0]music_select,
	 input rst_n,
	 output reg[511:0]row0,
	 output reg[511:0]row1,
	 output reg[511:0]row2,
	 output reg[511:0]row3,
	 output reg[511:0]row4,
	 output reg[511:0]row5,
	 output reg[511:0]row6,
	 output reg[511:0]row7,
	 output reg[511:0]row8,
	 output reg[511:0]row9,
	 output reg[511:0]row10,
	 output reg[511:0]row11,
	 output reg[511:0]row12,
	 output reg[511:0]row13,
	 output reg[511:0]row14,
	 output reg[511:0]row15,
	 output reg[511:0]row16,
	 output reg[511:0]row17,
	 output reg[511:0]row18,
	 output reg[511:0]row19,
	 output reg[511:0]row20,
	 output reg[511:0]row21,
	 output reg[511:0]row22,
	 output reg[511:0]row23,
	 output reg[511:0]row24,
	 output reg[511:0]row25,
	 output reg[511:0]row26,
	 output reg[511:0]row27,
	 output reg[511:0]row28,
	 output reg[511:0]row29,
	 output reg[511:0]row30,
	 output reg[511:0]row31,
	 output reg[511:0]row32,
	 output reg[511:0]row33,
	 output reg[511:0]row34,
	 output reg[511:0]row35,
	 output reg[511:0]row36,
	 output reg[511:0]row37,
	 output reg[511:0]row38,
	 output reg[511:0]row39,
	 output reg[511:0]row40,
	 output reg[511:0]row41,
	 output reg[511:0]row42,
	 output reg[511:0]row43,
	 output reg[511:0]row44,
	 output reg[511:0]row45,
	 output reg[511:0]row46,
	 output reg[511:0]row47,
	 output reg[511:0]row48,
	 output reg[511:0]row49,
	 output reg[511:0]row50,
	 output reg[511:0]row51,
	 output reg[511:0]row52,
	 output reg[511:0]row53,
	 output reg[511:0]row54,
	 output reg[511:0]row55,
	 output reg[511:0]row56,
	 output reg[511:0]row57,
	 output reg[511:0]row58,
	 output reg[511:0]row59,
	 output reg[511:0]row60,
	 output reg[511:0]row61,
	 output reg[511:0]row62,
	 output reg[511:0]row63
);
always@(*) begin
	if(!rst_n)begin
	row0<=0;
	row1<=0;
	row2<=0;
	row3<=0;
	row4<=0;
	row5<=0;
	row6<=0;
	row7<=0;
	row8<=0;
	row9<=0;
	row10<=0;
	row11<=0;
	row12<=0;
	row13<=0;
	row14<=0;
	row15<=0;
	row16<=0;
	row17<=0;
	row18<=0;
	row19<=0;
	row20<=0;
	row21<=0;
	row22<=0;
	row23<=0;
	row24<=0;
	row25<=0;
	row26<=0;
	row27<=0;
	row28<=0;
	row29<=0;
	row30<=0;
	row31<=0;
	row32<=0;
	row33<=0;
	row34<=0;
	row35<=0;
	row36<=0;
	row37<=0;
	row38<=0;
	row39<=0;
	row40<=0;
	row41<=0;
	row42<=0;
	row43<=0;
	row44<=0;
	row45<=0;
	row46<=0;
	row47<=0;
	row48<=0;
	row49<=0;
	row50<=0;
	row51<=0;
	row52<=0;
	row53<=0;
	row54<=0;
	row55<=0;
	row56<=0;
	row57<=0;
	row58<=0;
	row59<=0;
	row60<=0;
	row61<=0;
	row62<=0;
	row63<=0;
	end
	else begin
		case(music_select)
5'b00001:begin
row0<=512'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
row1<=512'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
row2<=512'h0000_0000_0000_0000_0000_0080_0400_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_4000_0800_0000_0000_0000;
row3<=512'h0000_0018_0000_0000_0000_00E0_0700_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0002_0000_0000_0000_E000_0E00_0000_0000_0000;
row4<=512'h0000_000E_0000_0000_0000_00F8_07C0_0000_0000_0000_0000_0000_0000_0000_0000_0800_0000_0003_8000_0000_0000_F800_0F00_0000_0000_0000;
row5<=512'h0000_0007_8000_0000_0000_00F0_07C0_0000_0000_0000_0000_0000_000C_0000_0000_1C00_0000_0003_F000_0000_0000_FC00_1FC0_0000_0000_0000;
row6<=512'h0000_0007_E000_0000_0000_00E0_0780_0000_0000_0000_0000_0000_000F_FFFF_FFFF_FF00_0000_0003_E000_0000_0001_F000_1F80_0000_0000_0000;
row7<=512'h0000_0003_E000_0000_0000_00E0_0780_0000_0000_0000_0000_0000_000F_FFFF_FFFF_FF00_0000_0003_C000_0000_0001_F000_1F00_0000_0000_0000;
row8<=512'h0000_0001_E000_0000_0000_00E0_0780_0000_0000_0000_0000_0000_000E_0000_0000_1E00_0000_0003_C000_0000_0001_E000_3F80_0000_0000_0000;
row9<=512'h0000_0001_E000_0000_0000_00E0_0780_0000_0000_0000_0000_0000_000E_0000_0000_1C00_0000_0003_C000_0000_0001_E000_3C80_0000_0000_0000;
row10<=512'h0000_0000_E000_0180_0000_00E0_0780_0000_0000_0000_0000_0000_000E_0001_C000_1C00_0000_0003_C000_0000_0003_C000_7CC0_0000_0000_0000;
row11<=512'h0000_0000_C000_07C0_0000_00E0_0780_0000_0000_0000_0000_0000_000E_0001_F000_1C00_0000_0003_C000_0400_0003_C000_7840_0000_0000_0000;
row12<=512'h0FFF_FFFF_FFFF_FFE0_0000_00E0_0780_0000_0000_0000_0000_0000_000E_0001_E000_1C00_0000_0003_C000_0E00_0003_8000_7860_0000_0000_0000;
row13<=512'h07FF_FFFF_FFFF_FFF0_0000_00E0_0780_0000_0000_0000_0000_0000_000E_0001_C000_1C00_0000_0003_C000_1F00_0007_8000_F030_0000_0000_0000;
row14<=512'h0200_3000_E000_0000_0000_00E0_0780_0800_0000_0000_0000_0000_000E_0001_C000_1C00_07FF_FFFF_FFFF_FF80_0007_0000_F030_0000_0000_0000;
row15<=512'h0000_3C00_F000_0000_0030_00E0_0780_1C00_0000_0000_0000_0000_000E_0001_C000_1C00_03FF_FFFF_FFFF_FFC0_000F_0001_E018_0000_0000_0000;
row16<=512'h0000_7E00_F800_0000_003F_FFFF_FFFF_FF00_0000_0000_0000_0000_000E_0001_C060_1C00_0100_001F_D000_0000_000F_0001_E01C_0000_0000_0000;
row17<=512'h0000_7C01_F000_0000_003F_FFFF_FFFF_FF00_0000_0000_0000_0000_000E_0001_C0F0_1C00_0000_001F_D800_0000_000E_0003_C00E_0000_0000_0000;
row18<=512'h0000_7801_E000_0000_003C_00E0_0780_1E00_0000_0000_0000_0000_000E_0FFF_FFF8_1C00_0000_003F_CC00_0000_001E_0003_800F_0000_0000_0000;
row19<=512'h0000_F801_E000_0000_003C_00E0_0780_1C00_0000_0000_0000_0000_000E_07FF_FFFC_1C00_0000_007F_CC00_0000_001C_0007_8007_8000_0000_0000;
row20<=512'h0000_F003_C000_2000_003C_00E0_0780_1C00_0000_0000_0000_0000_000E_0201_C000_1C00_0000_007B_C600_0000_003F_000F_0003_C000_0000_0000;
row21<=512'h0001_E003_C000_7000_003C_00E0_0780_1C00_0000_0000_0000_0000_000E_0001_C000_1C00_0000_00F3_C700_0000_003F_C00E_0003_E000_0000_0000;
row22<=512'h0001_E003_FFFF_FC00_003C_00E0_0780_1C00_0000_0000_0000_0000_000E_0001_C000_1C00_0000_01E3_C380_0000_0077_C01E_0001_F000_0000_0000;
row23<=512'h0001_C007_FFFF_FC00_003C_00E0_0780_1C00_0000_0000_0000_0000_000E_0001_C000_1C00_0000_03E3_C1C0_0000_0077_801C_0000_FC00_0000_0000;
row24<=512'h0003_C007_0000_7800_003C_00E0_0780_1C00_0000_0000_0000_0000_000E_0001_C000_1C00_0000_03C3_C1C0_0000_00E7_8038_0000_7E00_0000_0000;
row25<=512'h0003_800F_0000_F000_003C_00E0_0780_1C00_0000_0000_0000_0000_000E_0001_C00C_1C00_0000_0783_C0F0_0000_00C7_8070_0000_3F80_0000_0000;
row26<=512'h0007_800E_0000_F000_003C_00E0_0780_1C00_0000_0000_0000_0000_000E_0001_C01E_1C00_0000_0F03_C078_0000_01C7_80E0_0000_1FF0_0000_0000;
row27<=512'h0007_800E_3000_F000_003C_00E0_0780_1C00_0000_0000_0000_0000_000E_FFFF_FFFF_1C00_0000_1E03_C03C_0000_0187_80C4_0000_0FF8_0000_0000;
row28<=512'h000F_E01C_1801_E000_003C_00E0_0780_1C00_0000_0000_0000_0000_000E_7FFF_FFFF_9C00_0000_3C03_C03F_0000_0307_8187_0000_07C0_0000_0000;
row29<=512'h001F_E01C_1E01_E000_003C_00E0_0780_1C00_0000_0000_0000_0000_000E_3000_0000_1C00_0000_7803_C01F_8000_0707_8307_C000_0300_0000_0000;
row30<=512'h001F_C038_0F01_E000_003C_00E0_0780_1C00_0000_0000_0000_0000_000E_0000_0000_1C00_0000_F003_C00F_F000_0607_8607_C001_0000_0000_0000;
row31<=512'h003F_C03C_0783_C000_003C_00E0_0780_1C00_0000_0000_0000_0000_000E_0000_0000_1C00_0001_E003_C003_FC00_0C07_8C07_8003_8000_0000_0000;
row32<=512'h003B_C074_0783_C000_003C_00E0_0780_1C00_0000_0000_0000_0000_000E_0000_0000_1C00_0003_8003_C001_FFC0_1807_9807_8007_C000_0000_0000;
row33<=512'h0073_C0E6_0783_8000_003F_FFFF_FFFF_FC00_0000_0000_0000_0000_000E_0200_0040_1C00_000F_0003_C000_FFF8_1007_A007_800F_E000_0000_0000;
row34<=512'h00E3_C0E2_0387_8000_003F_FFFF_FFFF_FC00_0000_0000_0000_0000_000E_0180_00E0_1C00_001C_0003_C000_3FC0_0007_8007_801F_F000_0000_0000;
row35<=512'h00C3_C1C3_0387_8000_003C_00E0_0780_1C00_0000_0000_0000_0000_000E_01FF_FFF0_1C00_0038_0003_C000_0F80_0007_8007_803F_0000_0000_0000;
row36<=512'h01C3_C183_818F_0000_003C_00E0_0780_1C00_0000_0000_0000_0000_000E_01FF_FFF8_1C00_00E0_0003_C000_0300_0007_8007_807C_0000_0000_0000;
row37<=512'h0383_C301_810F_0000_003C_00E0_0780_1C00_0000_0000_0000_0000_001E_01C0_00E0_1C00_01C0_0003_C000_0000_0007_8007_81F0_0000_0000_0000;
row38<=512'h0303_C700_C01E_0000_003C_00E0_0780_1C00_0000_0000_0000_0000_001E_01C0_00E0_1C00_0700_0003_C000_0000_0007_8007_83C0_0000_0000_0000;
row39<=512'h0603_C600_E01E_0000_003C_00E0_0780_1C00_0000_0000_0000_0000_001C_01C0_00E0_1C00_1C00_0003_8000_0000_0007_8007_8F00_0000_0000_0000;
row40<=512'h0C03_CC00_603C_0000_003C_00E0_0780_1C00_0000_0000_0000_0000_001C_01C0_00E0_1C00_0000_0002_0000_0000_0007_8007_9C00_0000_0000_0000;
row41<=512'h0803_C800_703C_0000_003C_00E0_0780_1C00_0000_0000_0000_0000_001C_01C0_00E0_1C00_0000_0000_0000_0000_0007_8007_F000_0000_0000_0000;
row42<=512'h0003_C000_3878_0000_003C_00E0_0780_1C00_0000_0000_0000_0000_001C_01C0_00E0_1C00_0000_0000_0000_0000_0007_8007_C000_0000_0000_0000;
row43<=512'h0003_C000_3C78_0000_003C_00E0_0780_1C00_0000_0000_0000_0000_003C_01C0_00E0_1C00_0000_0000_0000_0000_0007_8007_8000_0000_0000_0000;
row44<=512'h0003_C000_1EF0_0000_003C_00E0_0780_1C00_0000_0000_0000_0000_0038_01C0_00E0_1C00_0004_0000_0001_0000_0007_8007_8000_0600_0000_0000;
row45<=512'h0003_C000_0FF0_0000_003C_00E0_0780_1C00_0000_0000_0000_0000_0038_01C0_00E0_1C00_0004_0200_1000_C000_0007_8007_8000_0600_0000_0000;
row46<=512'h0003_C000_0FE0_0000_003C_00E0_0780_1C00_0000_0000_0000_0000_0038_01FF_FFE0_1C00_000C_0300_1800_E000_0007_8007_8000_0600_0000_0000;
row47<=512'h0003_C000_07C0_0000_003C_00E0_0780_1C00_0000_0000_0000_0000_0070_01FF_FFE0_1C00_000C_0380_0E00_7000_0007_8007_8000_0600_0000_0000;
row48<=512'h0003_C000_07C0_0000_003C_00E0_0780_1C00_0000_0000_0000_0000_0070_01C0_00E0_1C00_000C_01C0_0F00_3800_0007_8007_8000_0600_0000_0000;
row49<=512'h0003_C000_0FF0_0000_003C_00E0_0780_1C00_0000_0000_0000_0000_0060_01C0_00E0_1C00_001C_01E0_0780_3E00_0007_8007_8000_0600_0000_0000;
row50<=512'h0003_C000_1FF8_0000_003C_00E0_0780_1C00_0000_0000_0000_0000_00E0_01C0_00F0_1C00_001C_00E0_07C0_1F00_0007_8007_8000_0600_0000_0000;
row51<=512'h0003_C000_3E7E_0000_003C_00E0_0780_1C00_0000_0000_0000_0000_00C0_01C0_0080_1C00_003C_00F0_03C0_1F00_0007_8007_8000_0600_0000_0000;
row52<=512'h0003_C000_7C3F_0000_003F_FFFF_FFFF_FC00_0000_0000_0000_0000_01C0_0100_0000_1C00_007C_00F8_03E0_0F80_0007_8007_8000_0E00_0000_0000;
row53<=512'h0003_C000_F01F_C000_003F_FFFF_FFFF_FC00_0000_0000_0000_0000_0180_0000_0000_1C00_0078_0078_03E0_0F80_0007_8007_8000_0E00_0000_0000;
row54<=512'h0003_C003_E00F_F800_003C_0000_0000_1C00_0000_0000_0000_0000_0380_0000_0000_3C00_00F8_0078_03E0_0780_0007_8007_8000_0F00_0000_0000;
row55<=512'h0003_C007_8003_FF80_003C_0000_0000_1C00_0000_0000_0000_0000_0300_0000_007F_FC00_01F8_0078_01C0_0780_0007_8007_C000_1FC0_0000_0000;
row56<=512'h0003_C01F_0001_FFF8_003C_0000_0000_1C00_0000_0000_0000_0000_0600_0000_000F_FC00_03F0_0070_0180_0780_0007_8003_FFFF_FF80_0000_0000;
row57<=512'h0003_C03C_0000_7FF0_003C_0000_0000_1C00_0000_0000_0000_0000_0600_0000_0003_F800_03E0_0060_0100_0300_0007_8003_FFFF_FF00_0000_0000;
row58<=512'h0003_C0F0_0000_1FC0_0038_0000_0000_1000_0000_0000_0000_0000_0C00_0000_0000_F000_0000_0000_0000_0200_0007_8000_FFFF_FE00_0000_0000;
row59<=512'h0003_C3C0_0000_0780_0020_0000_0000_0000_0000_0000_0000_0000_1800_0000_0000_E000_0000_0000_0000_0000_0007_8000_0000_0000_0000_0000;
row60<=512'h0003_8E00_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0007_0000_0000_0000_0000_0000;
row61<=512'h0002_1800_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0004_0000_0000_0000_0000_0000;
row62<=512'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
row63<=512'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
end
5'b00010:begin
row0<=512'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
row1<=512'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
row2<=512'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_4000_0800_0000_0000;
row3<=512'h0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0002_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0002_0000_0000_0000_E000_0E00_0000_0000;
row4<=512'h0000_001C_0000_0000_0000_0000_0000_0000_0000_0000_001F_0000_0000_0000_0000_0000_0000_0000_0000_0800_0000_0003_8000_0000_0000_F800_0F00_0000_0000;
row5<=512'h0000_001F_0000_0000_0004_0000_0000_8000_0000_0000_00FF_8000_0000_0000_0000_0000_000C_0000_0000_1C00_0000_0003_F000_0000_0000_FC00_1FC0_0000_0000;
row6<=512'h0000_001F_0000_0000_0002_0000_0001_C000_0000_0000_1FFF_E000_0000_0000_0000_0000_000F_FFFF_FFFF_FF00_0000_0003_E000_0000_0001_F000_1F80_0000_0000;
row7<=512'h0000_001E_0000_0000_0003_FFFF_FFFF_E000_0000_0007_FFFC_0000_0000_0000_0000_0000_000F_FFFF_FFFF_FF00_0000_0003_C000_0000_0001_F000_1F00_0000_0000;
row8<=512'h0000_001E_0000_0000_0003_FFFF_FFFF_F000_0000_03FF_FC00_0000_0000_0000_0000_0000_000E_0000_0000_1E00_0000_0003_C000_0000_0001_E000_3F80_0000_0000;
row9<=512'h0000_001E_0000_0000_0003_8003_8001_E000_0007_FFFF_C000_0000_0000_0000_0000_0000_000E_0000_0000_1C00_0000_0003_C000_0000_0001_E000_3C80_0000_0000;
row10<=512'h0000_001E_0000_0000_0003_8003_8001_C000_001C_0003_C000_0000_0000_0000_0000_0000_000E_0001_C000_1C00_0000_0003_C000_0000_0003_C000_7CC0_0000_0000;
row11<=512'h0000_001E_0000_0000_0003_8003_8001_C000_0000_0003_C000_0000_0000_0000_0000_0000_000E_0001_F000_1C00_0000_0003_C000_0400_0003_C000_7840_0000_0000;
row12<=512'h0000_001E_0000_0000_0003_8003_8001_C000_0000_0003_C000_0000_0000_0000_0000_0000_000E_0001_E000_1C00_0000_0003_C000_0E00_0003_8000_7860_0000_0000;
row13<=512'h0000_001E_0000_0000_0003_8003_8001_C000_0000_0003_C000_0000_0000_0000_0000_0000_000E_0001_C000_1C00_0000_0003_C000_1F00_0007_8000_F030_0000_0000;
row14<=512'h0000_001E_0000_0000_0003_8003_8001_C000_0000_0003_C000_0200_0000_0000_0000_0000_000E_0001_C000_1C00_07FF_FFFF_FFFF_FF80_0007_0000_F030_0000_0000;
row15<=512'h0000_001E_0000_0000_0003_8003_8001_C000_0000_0003_C000_0700_0000_0000_0000_0000_000E_0001_C000_1C00_03FF_FFFF_FFFF_FFC0_000F_0001_E018_0000_0000;
row16<=512'h0000_001E_0000_0000_0003_8003_8001_C000_0000_0003_C000_0F80_0000_0000_0000_0000_000E_0001_C060_1C00_0100_001F_D000_0000_000F_0001_E01C_0000_0000;
row17<=512'h0000_001E_0000_0600_0003_8003_8001_C000_0FFF_FFFF_FFFF_FFC0_0000_0000_0000_0000_000E_0001_C0F0_1C00_0000_001F_D800_0000_000E_0003_C00E_0000_0000;
row18<=512'h0000_001E_0000_0780_0003_8003_8001_C000_07FF_FFFF_FFFF_FFE0_0000_0000_0000_0000_000E_0FFF_FFF8_1C00_0000_003F_CC00_0000_001E_0003_800F_0000_0000;
row19<=512'h0000_001E_0000_0FE0_0003_FFFF_FFFF_C000_0200_003F_C800_0000_0000_0000_0000_0000_000E_07FF_FFFC_1C00_0000_007F_CC00_0000_001C_0007_8007_8000_0000;
row20<=512'h0000_001E_0000_1FE0_0003_FFFF_FFFF_C000_0000_007B_CC00_0000_0000_0000_0000_0000_000E_0201_C000_1C00_0000_007B_C600_0000_003F_000F_0003_C000_0000;
row21<=512'h0000_001E_0000_FE00_0003_8003_8001_C000_0000_00FB_C600_0000_0000_0000_0000_0000_000E_0001_C000_1C00_0000_00F3_C700_0000_003F_C00E_0003_E000_0000;
row22<=512'h0000_001E_000F_E000_0003_8003_8001_C000_0000_01F3_C700_0000_0000_0000_0000_0000_000E_0001_C000_1C00_0000_01E3_C380_0000_0077_C01E_0001_F000_0000;
row23<=512'h0000_001E_007E_0000_0003_8003_8001_C000_0000_03E3_C380_0000_0000_0000_0000_0000_000E_0001_C000_1C00_0000_03E3_C1C0_0000_0077_801C_0000_FC00_0000;
row24<=512'h0000_001E_07E0_0000_0003_8003_8001_C000_0000_07C3_C1C0_0000_0000_0000_0000_0000_000E_0001_C000_1C00_0000_03C3_C1C0_0000_00E7_8038_0000_7E00_0000;
row25<=512'h0000_001E_7E00_0000_0003_8003_8001_C000_0000_0F03_C0F0_0000_0000_0000_0000_0000_000E_0001_C00C_1C00_0000_0783_C0F0_0000_00C7_8070_0000_3F80_0000;
row26<=512'h0000_001F_E000_0000_0003_8003_8001_C000_0000_1E03_C078_0000_0000_0000_0000_0000_000E_0001_C01E_1C00_0000_0F03_C078_0000_01C7_80E0_0000_1FF0_0000;
row27<=512'h0000_007E_0000_0000_0003_8003_8001_C000_0000_3C03_C03E_0000_0000_0000_0000_0000_000E_FFFF_FFFF_1C00_0000_1E03_C03C_0000_0187_80C4_0000_0FF8_0000;
row28<=512'h0000_07FE_0000_0000_0003_8003_8001_C000_0000_7803_C01F_8000_0000_0000_0000_0000_000E_7FFF_FFFF_9C00_0000_3C03_C03F_0000_0307_8187_0000_07C0_0000;
row29<=512'h0000_7E1E_0000_0000_0003_8003_8001_C000_0001_F003_C00F_F000_0000_0000_0000_0000_000E_3000_0000_1C00_0000_7803_C01F_8000_0707_8307_C000_0300_0000;
row30<=512'h0007_E01E_0000_0000_0003_8003_8001_C000_0003_C003_C003_FE00_0000_0000_0000_0000_000E_0000_0000_1C00_0000_F003_C00F_F000_0607_8607_C001_0000_0000;
row31<=512'h00FE_001E_0000_0000_0003_8003_8001_C000_0007_8003_C001_FFE0_0000_0000_0000_0000_000E_0000_0000_1C00_0001_E003_C003_FC00_0C07_8C07_8003_8000_0000;
row32<=512'h0FE0_001E_0000_0000_0003_FFFF_FFFF_C000_001E_0003_0000_7FF8_0000_0000_0000_0000_000E_0000_0000_1C00_0003_8003_C001_FFC0_1807_9807_8007_C000_0000;
row33<=512'h1F00_001E_0000_0000_0003_FFFF_FFFF_C000_0038_0000_000C_1FC0_0000_0000_0000_0000_000E_0200_0040_1C00_000F_0003_C000_FFF8_1007_A007_800F_E000_0000;
row34<=512'h0400_001E_0000_0000_0003_8003_8001_C000_00F0_6000_000E_0780_0000_0000_0000_0000_000E_0180_00E0_1C00_001C_0003_C000_3FC0_0007_8007_801F_F000_0000;
row35<=512'h0000_001E_0000_0000_0003_8003_8001_C000_01C0_7FFF_FFFF_0100_0000_0000_0000_0000_000E_01FF_FFF0_1C00_0038_0003_C000_0F80_0007_8007_803F_0000_0000;
row36<=512'h0000_001E_0000_0000_0003_8003_8001_8000_0700_7FFF_FFFF_0000_0000_0000_0000_0000_000E_01FF_FFF8_1C00_00E0_0003_C000_0300_0007_8007_807C_0000_0000;
row37<=512'h0000_001E_0000_0000_0002_0003_8000_0000_1C00_7800_001E_0000_0000_0000_0000_0000_001E_01C0_00E0_1C00_01C0_0003_C000_0000_0007_8007_81F0_0000_0000;
row38<=512'h0000_001E_0000_0000_0000_0003_8000_0000_1000_7800_001E_0000_0000_0000_0000_0000_001E_01C0_00E0_1C00_0700_0003_C000_0000_0007_8007_83C0_0000_0000;
row39<=512'h0000_001E_0000_0080_0000_0003_8000_0000_0000_7800_001E_0000_0000_0000_0000_0000_001C_01C0_00E0_1C00_1C00_0003_8000_0000_0007_8007_8F00_0000_0000;
row40<=512'h0000_001E_0000_0080_0000_0003_8000_0000_0000_7800_001E_0000_0000_0000_0000_0000_001C_01C0_00E0_1C00_0000_0002_0000_0000_0007_8007_9C00_0000_0000;
row41<=512'h0000_001E_0000_0080_0000_0003_8000_2000_0000_7800_001E_0000_0000_0000_0000_0000_001C_01C0_00E0_1C00_0000_0000_0000_0000_0007_8007_F000_0000_0000;
row42<=512'h0000_001E_0000_0080_0000_0003_8000_7000_0000_7800_001E_0000_0000_0000_0000_0000_001C_01C0_00E0_1C00_0000_0000_0000_0000_0007_8007_C000_0000_0000;
row43<=512'h0000_001E_0000_0080_0000_0003_8000_F800_0000_7800_001E_0000_0000_0000_0000_0000_003C_01C0_00E0_1C00_0000_0000_0000_0000_0007_8007_8000_0000_0000;
row44<=512'h0000_001E_0000_00C0_007F_FFFF_FFFF_FC00_0000_7800_001E_0000_0000_0000_0000_0000_0038_01C0_00E0_1C00_0004_0000_0001_0000_0007_8007_8000_0600_0000;
row45<=512'h0000_001E_0000_00C0_003F_FFFF_FFFF_FE00_0000_7FFF_FFFE_0000_0000_0000_0000_0000_0038_01C0_00E0_1C00_0004_0200_1000_C000_0007_8007_8000_0600_0000;
row46<=512'h0000_001E_0000_01C0_0010_0003_8000_0000_0000_7FFF_FFFE_0000_0000_0000_0000_0000_0038_01FF_FFE0_1C00_000C_0300_1800_E000_0007_8007_8000_0600_0000;
row47<=512'h0000_001E_0000_01C0_0000_0003_8000_0000_0000_7800_001E_0000_0000_0000_0000_0000_0070_01FF_FFE0_1C00_000C_0380_0E00_7000_0007_8007_8000_0600_0000;
row48<=512'h0000_001E_0000_01C0_0000_0003_8000_0000_0000_7800_001E_0000_0000_0000_0000_0000_0070_01C0_00E0_1C00_000C_01C0_0F00_3800_0007_8007_8000_0600_0000;
row49<=512'h0000_001E_0000_01C0_0000_0003_8000_0000_0000_7800_001E_0000_0000_0000_0000_0000_0060_01C0_00E0_1C00_001C_01E0_0780_3E00_0007_8007_8000_0600_0000;
row50<=512'h0000_001E_0000_01C0_0000_0003_8000_0000_0000_7800_001E_0000_0000_0000_0000_0000_00E0_01C0_00F0_1C00_001C_00E0_07C0_1F00_0007_8007_8000_0600_0000;
row51<=512'h0000_001E_0000_01E0_0000_0003_8000_0000_0000_7800_001E_0000_0000_0000_0000_0000_00C0_01C0_0080_1C00_003C_00F0_03C0_1F00_0007_8007_8000_0600_0000;
row52<=512'h0000_001F_0000_03F0_0000_0003_8000_0000_0000_7800_001E_0000_0000_0000_0000_0000_01C0_0100_0000_1C00_007C_00F8_03E0_0F80_0007_8007_8000_0E00_0000;
row53<=512'h0000_001F_8000_07F8_0000_0003_8000_0000_0000_7800_001E_0000_0000_0000_0000_0000_0180_0000_0000_1C00_0078_0078_03E0_0F80_0007_8007_8000_0E00_0000;
row54<=512'h0000_000F_FFFF_FFF8_0000_0003_8000_0180_0000_7FFF_FFFE_0000_0000_0000_0000_0000_0380_0000_0000_3C00_00F8_0078_03E0_0780_0007_8007_8000_0F00_0000;
row55<=512'h0000_0007_FFFF_FFF0_0000_0003_8000_03C0_0000_7FFF_FFFE_0000_0000_0000_0000_0000_0300_0000_007F_FC00_01F8_0078_01C0_0780_0007_8007_C000_1FC0_0000;
row56<=512'h0000_0001_FFFF_FF80_0000_0003_8000_07E0_0000_7800_001E_0000_0000_0000_0000_0000_0600_0000_000F_FC00_03F0_0070_0180_0780_0007_8003_FFFF_FF80_0000;
row57<=512'h0000_0000_0000_0000_1FFF_FFFF_FFFF_FFF0_0000_7800_001E_0000_0000_0000_0000_0000_0600_0000_0003_F800_03E0_0060_0100_0300_0007_8003_FFFF_FF00_0000;
row58<=512'h0000_0000_0000_0000_0FFF_FFFF_FFFF_FFF8_0000_7800_001E_0000_0000_0000_0000_0000_0C00_0000_0000_F000_0000_0000_0000_0200_0007_8000_FFFF_FE00_0000;
row59<=512'h0000_0000_0000_0000_0600_0000_0000_0000_0000_7000_001C_0000_0000_0000_0000_0000_1800_0000_0000_E000_0000_0000_0000_0000_0007_8000_0000_0000_0000;
row60<=512'h0000_0000_0000_0000_0000_0000_0000_0000_0000_4000_0010_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0007_0000_0000_0000_0000;
row61<=512'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0004_0000_0000_0000_0000;
row62<=512'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
row63<=512'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
end
5'b00100:begin
row0<=512'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
row1<=512'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
row2<=512'h0000_0008_0000_0000_0000_0000_0200_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_4000_0800_0000_0000_0000;
row3<=512'h0000_0006_0000_0000_0000_C000_0300_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0002_0000_0000_0000_E000_0E00_0000_0000_0000;
row4<=512'h0000_0007_0000_0000_0000_F000_07C0_0000_0000_0000_0000_0000_0000_0000_0000_0800_0000_0003_8000_0000_0000_F800_0F00_0000_0000_0000;
row5<=512'h0000_0003_C000_0000_0000_F000_07C0_0000_0000_0000_0000_0000_000C_0000_0000_1C00_0000_0003_F000_0000_0000_FC00_1FC0_0000_0000_0000;
row6<=512'h0000_0001_E000_0000_0000_E000_0780_0000_0000_0000_0000_0000_000F_FFFF_FFFF_FF00_0000_0003_E000_0000_0001_F000_1F80_0000_0000_0000;
row7<=512'h0000_0001_E000_0000_0000_E000_0F00_0000_0000_0000_0000_0000_000F_FFFF_FFFF_FF00_0000_0003_C000_0000_0001_F000_1F00_0000_0000_0000;
row8<=512'h0000_0000_F000_0000_0000_E010_0E00_4000_0000_0000_0000_0000_000E_0000_0000_1E00_0000_0003_C000_0000_0001_E000_3F80_0000_0000_0000;
row9<=512'h0000_0000_F000_0000_0000_E038_1E00_E000_0000_0000_0000_0000_000E_0000_0000_1C00_0000_0003_C000_0000_0001_E000_3C80_0000_0000_0000;
row10<=512'h0004_0000_F000_0000_0FFF_FFFC_1FFF_F000_0000_0000_0000_0000_000E_0001_C000_1C00_0000_0003_C000_0000_0003_C000_7CC0_0000_0000_0000;
row11<=512'h0004_0000_E000_0600_07FF_FFFE_3FFF_F800_0000_0000_0000_0000_000E_0001_F000_1C00_0000_0003_C000_0400_0003_C000_7840_0000_0000_0000;
row12<=512'h000C_0000_4000_0F00_0300_E000_3801_F000_0000_0000_0000_0000_000E_0001_E000_1C00_0000_0003_C000_0E00_0003_8000_7860_0000_0000_0000;
row13<=512'h000F_FFFF_FFFF_FF80_0000_E000_7001_C000_0000_0000_0000_0000_000E_0001_C000_1C00_0000_0003_C000_1F00_0007_8000_F030_0000_0000_0000;
row14<=512'h000F_FFFF_FFFF_FFC0_0000_E000_7003_8000_0000_0000_0000_0000_000E_0001_C000_1C00_07FF_FFFF_FFFF_FF80_0007_0000_F030_0000_0000_0000;
row15<=512'h001C_0000_0000_0F80_0000_E000_E003_0000_0000_0000_0000_0000_000E_0001_C000_1C00_03FF_FFFF_FFFF_FFC0_000F_0001_E018_0000_0000_0000;
row16<=512'h001C_0000_0000_1E00_0000_E060_C006_0000_0000_0000_0000_0000_000E_0001_C060_1C00_0100_001F_D000_0000_000F_0001_E01C_0000_0000_0000;
row17<=512'h003C_0000_0000_1C00_03FF_FFF1_8006_0000_0000_0000_0000_0000_000E_0001_C0F0_1C00_0000_001F_D800_0000_000E_0003_C00E_0000_0000_0000;
row18<=512'h007C_0000_0000_1800_01FF_FFFB_000C_0400_0000_0000_0000_0000_000E_0FFF_FFF8_1C00_0000_003F_CC00_0000_001E_0003_800F_0000_0000_0000;
row19<=512'h00FC_0020_0000_3000_0080_E006_0008_0E00_0000_0000_0000_0000_000E_07FF_FFFC_1C00_0000_007F_CC00_0000_001C_0007_8007_8000_0000_0000;
row20<=512'h01F8_0038_0000_2000_0000_E005_FFFF_FF00_0000_0000_0000_0000_000E_0201_C000_1C00_0000_007B_C600_0000_003F_000F_0003_C000_0000_0000;
row21<=512'h0070_003E_0000_4000_0000_E000_FFFF_FF80_0000_0000_0000_0000_000E_0001_C000_1C00_0000_00F3_C700_0000_003F_C00E_0003_E000_0000_0000;
row22<=512'h0000_003E_0000_0000_0000_E008_6070_0F00_0000_0000_0000_0000_000E_0001_C000_1C00_0000_01E3_C380_0000_0077_C01E_0001_F000_0000_0000;
row23<=512'h0000_007C_0000_0000_0000_E01C_0070_0E00_0000_0000_0000_0000_000E_0001_C000_1C00_0000_03E3_C1C0_0000_0077_801C_0000_FC00_0000_0000;
row24<=512'h0000_0078_0000_0000_1FFF_FFFE_0070_0E00_0000_0000_0000_0000_000E_0001_C000_1C00_0000_03C3_C1C0_0000_00E7_8038_0000_7E00_0000_0000;
row25<=512'h0000_0078_0000_0000_0FFF_FFFF_0070_0E00_0000_0000_0000_0000_000E_0001_C00C_1C00_0000_0783_C0F0_0000_00C7_8070_0000_3F80_0000_0000;
row26<=512'h0000_00F0_0000_0300_0400_0000_0070_0E00_0000_0000_0000_0000_000E_0001_C01E_1C00_0000_0F03_C078_0000_01C7_80E0_0000_1FF0_0000_0000;
row27<=512'h0000_00F0_0000_0780_0000_0000_0070_0E00_0000_0000_0000_0000_000E_FFFF_FFFF_1C00_0000_1E03_C03C_0000_0187_80C4_0000_0FF8_0000_0000;
row28<=512'h0000_00E0_0000_0FC0_0100_0040_0070_0E40_0000_0000_0000_0000_000E_7FFF_FFFF_9C00_0000_3C03_C03F_0000_0307_8187_0000_07C0_0000_0000;
row29<=512'h0FFF_FFFF_FFFF_FFE0_0180_00E0_0070_0EE0_0000_0000_0000_0000_000E_3000_0000_1C00_0000_7803_C01F_8000_0707_8307_C000_0300_0000_0000;
row30<=512'h07FF_FFFF_FFFF_FFF0_01FF_FFF7_FFFF_FFF0_0000_0000_0000_0000_000E_0000_0000_1C00_0000_F003_C00F_F000_0607_8607_C001_0000_0000_0000;
row31<=512'h0000_01C0_003E_0000_01FF_FFFB_FFFF_FFF8_0000_0000_0000_0000_000E_0000_0000_1C00_0001_E003_C003_FC00_0C07_8C07_8003_8000_0000_0000;
row32<=512'h0000_03C0_003C_0000_01E0_01E1_0070_0E00_0000_0000_0000_0000_000E_0000_0000_1C00_0003_8003_C001_FFC0_1807_9807_8007_C000_0000_0000;
row33<=512'h0000_0380_007C_0000_01E0_01E0_0070_0E00_0000_0000_0000_0000_000E_0200_0040_1C00_000F_0003_C000_FFF8_1007_A007_800F_E000_0000_0000;
row34<=512'h0000_0780_0078_0000_01E0_01E0_0070_0E00_0000_0000_0000_0000_000E_0180_00E0_1C00_001C_0003_C000_3FC0_0007_8007_801F_F000_0000_0000;
row35<=512'h0000_0700_00F8_0000_01E0_01E0_0070_0E00_0000_0000_0000_0000_000E_01FF_FFF0_1C00_0038_0003_C000_0F80_0007_8007_803F_0000_0000_0000;
row36<=512'h0000_0F00_00F0_0000_01E0_01E0_0070_0E00_0000_0000_0000_0000_000E_01FF_FFF8_1C00_00E0_0003_C000_0300_0007_8007_807C_0000_0000_0000;
row37<=512'h0000_0E00_01F0_0000_01FF_FFE0_0070_0E00_0000_0000_0000_0000_001E_01C0_00E0_1C00_01C0_0003_C000_0000_0007_8007_81F0_0000_0000_0000;
row38<=512'h0000_1E00_01E0_0000_01FF_FFE0_0070_0E00_0000_0000_0000_0000_001E_01C0_00E0_1C00_0700_0003_C000_0000_0007_8007_83C0_0000_0000_0000;
row39<=512'h0000_1C00_03E0_0000_01E0_01E0_0070_0E00_0000_0000_0000_0000_001C_01C0_00E0_1C00_1C00_0003_8000_0000_0007_8007_8F00_0000_0000_0000;
row40<=512'h0000_3C00_03C0_0000_01E0_01E0_0070_0E00_0000_0000_0000_0000_001C_01C0_00E0_1C00_0000_0002_0000_0000_0007_8007_9C00_0000_0000_0000;
row41<=512'h0000_3800_0780_0000_01E0_01E3_FFFF_FE00_0000_0000_0000_0000_001C_01C0_00E0_1C00_0000_0000_0000_0000_0007_8007_F000_0000_0000_0000;
row42<=512'h0000_7800_0780_0000_01E0_01E1_FFFF_FE00_0000_0000_0000_0000_001C_01C0_00E0_1C00_0000_0000_0000_0000_0007_8007_C000_0000_0000_0000;
row43<=512'h0000_7F80_0F00_0000_01E0_01E0_C070_0E00_0000_0000_0000_0000_003C_01C0_00E0_1C00_0000_0000_0000_0000_0007_8007_8000_0000_0000_0000;
row44<=512'h0000_03FC_1F00_0000_01E0_01E0_0070_0C00_0000_0000_0000_0000_0038_01C0_00E0_1C00_0004_0000_0001_0000_0007_8007_8000_0600_0000_0000;
row45<=512'h0000_007F_BE00_0000_01FF_FFE0_0070_0000_0000_0000_0000_0000_0038_01C0_00E0_1C00_0004_0200_1000_C000_0007_8007_8000_0600_0000_0000;
row46<=512'h0000_0007_FC00_0000_01FF_FFE0_0070_0000_0000_0000_0000_0000_0038_01FF_FFE0_1C00_000C_0300_1800_E000_0007_8007_8000_0600_0000_0000;
row47<=512'h0000_0000_FF00_0000_01E0_01E0_0070_0000_0000_0000_0000_0000_0070_01FF_FFE0_1C00_000C_0380_0E00_7000_0007_8007_8000_0600_0000_0000;
row48<=512'h0000_0000_FFE0_0000_01E0_01E0_0070_0000_0000_0000_0000_0000_0070_01C0_00E0_1C00_000C_01C0_0F00_3800_0007_8007_8000_0600_0000_0000;
row49<=512'h0000_0001_F7FC_0000_01E0_01E0_0070_0000_0000_0000_0000_0000_0060_01C0_00E0_1C00_001C_01E0_0780_3E00_0007_8007_8000_0600_0000_0000;
row50<=512'h0000_0003_E1FF_0000_01E0_01E0_0070_0000_0000_0000_0000_0000_00E0_01C0_00F0_1C00_001C_00E0_07C0_1F00_0007_8007_8000_0600_0000_0000;
row51<=512'h0000_0007_C03F_C000_01E0_01E0_0070_0000_0000_0000_0000_0000_00C0_01C0_0080_1C00_003C_00F0_03C0_1F00_0007_8007_8000_0600_0000_0000;
row52<=512'h0000_001F_000F_F800_01E0_01E0_0070_0000_0000_0000_0000_0000_01C0_0100_0000_1C00_007C_00F8_03E0_0F80_0007_8007_8000_0E00_0000_0000;
row53<=512'h0000_007E_0003_FC00_01E0_01E0_0070_0000_0000_0000_0000_0000_0180_0000_0000_1C00_0078_0078_03E0_0F80_0007_8007_8000_0E00_0000_0000;
row54<=512'h0000_01F8_0001_FE00_01E0_01E0_0070_0000_0000_0000_0000_0000_0380_0000_0000_3C00_00F8_0078_03E0_0780_0007_8007_8000_0F00_0000_0000;
row55<=512'h0000_07E0_0000_7F00_01E0_01E0_0070_0000_0000_0000_0000_0000_0300_0000_007F_FC00_01F8_0078_01C0_0780_0007_8007_C000_1FC0_0000_0000;
row56<=512'h0000_1F80_0000_3F80_01E0_E1C0_F0F0_0000_0000_0000_0000_0000_0600_0000_000F_FC00_03F0_0070_0180_0780_0007_8003_FFFF_FF80_0000_0000;
row57<=512'h0000_FE00_0000_1F80_01E0_7FC0_3FF0_0000_0000_0000_0000_0000_0600_0000_0003_F800_03E0_0060_0100_0300_0007_8003_FFFF_FF00_0000_0000;
row58<=512'h000F_E000_0000_0780_01E0_1FC0_0FF0_0000_0000_0000_0000_0000_0C00_0000_0000_F000_0000_0000_0000_0200_0007_8000_FFFF_FE00_0000_0000;
row59<=512'h00FF_0000_0000_0100_01E0_0F80_07E0_0000_0000_0000_0000_0000_1800_0000_0000_E000_0000_0000_0000_0000_0007_8000_0000_0000_0000_0000;
row60<=512'h07C0_0000_0000_0000_0180_0700_03C0_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0007_0000_0000_0000_0000_0000;
row61<=512'h0000_0000_0000_0000_0100_0400_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0004_0000_0000_0000_0000_0000;
row62<=512'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
row63<=512'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
end
5'b01000:begin
row0<=512'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
row1<=512'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
row2<=512'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_4000_0800_0000_0000_0000;
row3<=512'h0002_0000_0000_0000_0000_0000_3000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0002_0000_0000_0000_E000_0E00_0000_0000_0000;
row4<=512'h0003_8000_0700_0000_0180_0000_1C00_0000_0000_0000_0000_0000_0000_0000_0000_0800_0000_0003_8000_0000_0000_F800_0F00_0000_0000_0000;
row5<=512'h0007_C000_07C0_0000_00E0_0000_0E00_0000_0000_0000_0000_0000_000C_0000_0000_1C00_0000_0003_F000_0000_0000_FC00_1FC0_0000_0000_0000;
row6<=512'h0007_E000_07C0_0000_0078_0000_0F80_0000_0000_0000_0000_0000_000F_FFFF_FFFF_FF00_0000_0003_E000_0000_0001_F000_1F80_0000_0000_0000;
row7<=512'h0007_8000_0780_0000_003C_0000_07C0_0000_0000_0000_0000_0000_000F_FFFF_FFFF_FF00_0000_0003_C000_0000_0001_F000_1F00_0000_0000_0000;
row8<=512'h0007_8000_0700_0000_003E_0000_07C0_0000_0000_0000_0000_0000_000E_0000_0000_1E00_0000_0003_C000_0000_0001_E000_3F80_0000_0000_0000;
row9<=512'h0007_0000_0700_0000_001F_0000_03C0_0000_0000_0000_0000_0000_000E_0000_0000_1C00_0000_0003_C000_0000_0001_E000_3C80_0000_0000_0000;
row10<=512'h000F_0000_0700_0000_001F_0000_03C0_0000_0000_0000_0000_0000_000E_0001_C000_1C00_0000_0003_C000_0000_0003_C000_7CC0_0000_0000_0000;
row11<=512'h000F_0000_0700_0000_000F_0000_01C0_0080_0000_0000_0000_0000_000E_0001_F000_1C00_0000_0003_C000_0400_0003_C000_7840_0000_0000_0000;
row12<=512'h000E_0030_0700_0000_000F_0000_01C0_01C0_0000_0000_0000_0000_000E_0001_E000_1C00_0000_0003_C000_0E00_0003_8000_7860_0000_0000_0000;
row13<=512'h000E_0078_0700_0000_000E_1FFF_FFFF_FFE0_0000_0000_0000_0000_000E_0001_C000_1C00_0000_0003_C000_1F00_0007_8000_F030_0000_0000_0000;
row14<=512'h1FFF_FFFC_0700_0000_0004_0FFF_FFFF_FFF0_0000_0000_0000_0000_000E_0001_C000_1C00_07FF_FFFF_FFFF_FF80_0007_0000_F030_0000_0000_0000;
row15<=512'h0FFF_FFFE_0700_0000_0000_0600_F00F_0000_0000_0000_0000_0000_000E_0001_C000_1C00_03FF_FFFF_FFFF_FFC0_000F_0001_E018_0000_0000_0000;
row16<=512'h041C_0000_0700_C000_0000_0000_F00F_0000_0000_0000_0000_0000_000E_0001_C060_1C00_0100_001F_D000_0000_000F_0001_E01C_0000_0000_0000;
row17<=512'h003C_0000_0700_E000_0000_0000_F00F_0000_0000_0000_0000_0000_000E_0001_C0F0_1C00_0000_001F_D800_0000_000E_0003_C00E_0000_0000_0000;
row18<=512'h003C_0000_0701_F800_0000_0000_F00F_0000_0000_0000_0000_0000_000E_0FFF_FFF8_1C00_0000_003F_CC00_0000_001E_0003_800F_0000_0000_0000;
row19<=512'h0038_4000_3FFF_F000_0000_0000_F00F_0000_0000_0000_0000_0000_000E_07FF_FFFC_1C00_0000_007F_CC00_0000_001C_0007_8007_8000_0000_0000;
row20<=512'h0078_700F_FF01_E000_0000_0000_F00F_0000_0000_0000_0000_0000_000E_0201_C000_1C00_0000_007B_C600_0000_003F_000F_0003_C000_0000_0000;
row21<=512'h0078_7C02_0701_C000_0000_0040_F00F_0000_0000_0000_0000_0000_000E_0001_C000_1C00_0000_00F3_C700_0000_003F_C00E_0003_E000_0000_0000;
row22<=512'h0070_7C00_0701_C000_0002_0070_F00F_0000_0000_0000_0000_0000_000E_0001_C000_1C00_0000_01E3_C380_0000_0077_C01E_0001_F000_0000_0000;
row23<=512'h00F0_7000_0701_C000_0007_007C_F00F_4000_0000_0000_0000_0000_000E_0001_C000_1C00_0000_03E3_C1C0_0000_0077_801C_0000_FC00_0000_0000;
row24<=512'h00F0_7000_0701_C000_3FFF_807C_F00F_3000_0000_0000_0000_0000_000E_0001_C000_1C00_0000_03C3_C1C0_0000_00E7_8038_0000_7E00_0000_0000;
row25<=512'h00E0_7000_0701_C000_1FFF_C0F0_F00F_1800_0000_0000_0000_0000_000E_0001_C00C_1C00_0000_0783_C0F0_0000_00C7_8070_0000_3F80_0000_0000;
row26<=512'h01E0_7000_0701_C000_0C0F_80F0_F00F_1C00_0000_0000_0000_0000_000E_0001_C01E_1C00_0000_0F03_C078_0000_01C7_80E0_0000_1FF0_0000_0000;
row27<=512'h03C0_7020_0701_C000_000F_01E0_F00F_0E00_0000_0000_0000_0000_000E_FFFF_FFFF_1C00_0000_1E03_C03C_0000_0187_80C4_0000_0FF8_0000_0000;
row28<=512'h03C0_7070_0701_C000_000F_01C0_F00F_0700_0000_0000_0000_0000_000E_7FFF_FFFF_9C00_0000_3C03_C03F_0000_0307_8187_0000_07C0_0000_0000;
row29<=512'h0FFF_FFF8_0701_C000_000F_01C0_F00F_0780_0000_0000_0000_0000_000E_3000_0000_1C00_0000_7803_C01F_8000_0707_8307_C000_0300_0000_0000;
row30<=512'h07FF_FFFC_0F01_C000_000F_0380_F00F_03C0_0000_0000_0000_0000_000E_0000_0000_1C00_0000_F003_C00F_F000_0607_8607_C001_0000_0000_0000;
row31<=512'h0380_7000_0F01_C000_000F_0300_E00F_03E0_0000_0000_0000_0000_000E_0000_0000_1C00_0001_E003_C003_FC00_0C07_8C07_8003_8000_0000_0000;
row32<=512'h0100_7000_0E01_C000_000F_0700_E00F_01E0_0000_0000_0000_0000_000E_0000_0000_1C00_0003_8003_C001_FFC0_1807_9807_8007_C000_0000_0000;
row33<=512'h0000_7000_0E01_C000_000F_0E00_E00F_01E0_0000_0000_0000_0000_000E_0200_0040_1C00_000F_0003_C000_FFF8_1007_A007_800F_E000_0000_0000;
row34<=512'h0000_7000_0E01_C000_000F_0C01_E00F_00E0_0000_0000_0000_0000_000E_0180_00E0_1C00_001C_0003_C000_3FC0_0007_8007_801F_F000_0000_0000;
row35<=512'h0000_7000_0E01_C000_000F_1801_E00F_00E0_0000_0000_0000_0000_000E_01FF_FFF0_1C00_0038_0003_C000_0F80_0007_8007_803F_0000_0000_0000;
row36<=512'h0000_7000_1E01_C000_000F_3001_C00F_00C0_0000_0000_0000_0000_000E_01FF_FFF8_1C00_00E0_0003_C000_0300_0007_8007_807C_0000_0000_0000;
row37<=512'h0000_7000_1C01_C000_000F_2003_C00F_0000_0000_0000_0000_0000_001E_01C0_00E0_1C00_01C0_0003_C000_0000_0007_8007_81F0_0000_0000_0000;
row38<=512'h0000_7004_1C01_C000_000F_0003_800F_0000_0000_0000_0000_0000_001E_01C0_00E0_1C00_0700_0003_C000_0000_0007_8007_83C0_0000_0000_0000;
row39<=512'h0000_707C_1C01_C000_000F_0003_800F_0000_0000_0000_0000_0000_001C_01C0_00E0_1C00_1C00_0003_8000_0000_0007_8007_8F00_0000_0000_0000;
row40<=512'h0000_73E0_3C01_C000_000F_0007_000F_0000_0000_0000_0000_0000_001C_01C0_00E0_1C00_0000_0002_0000_0000_0007_8007_9C00_0000_0000_0000;
row41<=512'h0000_7F80_3801_C000_000F_000F_000F_0000_0000_0000_0000_0000_001C_01C0_00E0_1C00_0000_0000_0000_0000_0007_8007_F000_0000_0000_0000;
row42<=512'h0003_FC00_3801_C000_000F_000E_000F_0000_0000_0000_0000_0000_001C_01C0_00E0_1C00_0000_0000_0000_0000_0007_8007_C000_0000_0000_0000;
row43<=512'h003F_F000_7001_C000_000F_001C_000F_0000_0000_0000_0000_0000_003C_01C0_00E0_1C00_0000_0000_0000_0000_0007_8007_8000_0000_0000_0000;
row44<=512'h03FF_7000_7001_C000_000F_0038_000F_0000_0000_0000_0000_0000_0038_01C0_00E0_1C00_0004_0000_0001_0000_0007_8007_8000_0600_0000_0000;
row45<=512'h0FFC_7000_F001_C040_000F_0070_000F_0000_0000_0000_0000_0000_0038_01C0_00E0_1C00_0004_0200_1000_C000_0007_8007_8000_0600_0000_0000;
row46<=512'h0FF0_7000_E001_C040_000F_00E0_1F1F_0000_0000_0000_0000_0000_0038_01FF_FFE0_1C00_000C_0300_1800_E000_0007_8007_8000_0600_0000_0000;
row47<=512'h07C0_7000_E001_C040_000F_01C0_03FE_0000_0000_0000_0000_0000_0070_01FF_FFE0_1C00_000C_0380_0E00_7000_0007_8007_8000_0600_0000_0000;
row48<=512'h0700_7001_C001_C040_001F_8300_00FE_0000_0000_0000_0000_0000_0070_01C0_00E0_1C00_000C_01C0_0F00_3800_0007_8007_8000_0600_0000_0000;
row49<=512'h0000_7003_8001_C060_0078_E600_007E_0000_0000_0000_0000_0000_0060_01C0_00E0_1C00_001C_01E0_0780_3E00_0007_8007_8000_0600_0000_0000;
row50<=512'h0000_7003_8001_C060_00F0_7000_003C_0000_0000_0000_0000_0000_00E0_01C0_00F0_1C00_001C_00E0_07C0_1F00_0007_8007_8000_0600_0000_0000;
row51<=512'h0000_7007_0001_C060_03E0_1C00_0018_0000_0000_0000_0000_0000_00C0_01C0_0080_1C00_003C_00F0_03C0_1F00_0007_8007_8000_0600_0000_0000;
row52<=512'h0000_7006_0001_C060_07C0_0F80_0000_0000_0000_0000_0000_0000_01C0_0100_0000_1C00_007C_00F8_03E0_0F80_0007_8007_8000_0E00_0000_0000;
row53<=512'h0000_700C_0001_E0F0_1F80_03F8_0000_007C_0000_0000_0000_0000_0180_0000_0000_1C00_0078_0078_03E0_0F80_0007_8007_8000_0E00_0000_0000;
row54<=512'h0000_701C_0001_FFF8_1F00_01FF_FFFF_FFF0_0000_0000_0000_0000_0380_0000_0000_3C00_00F8_0078_03E0_0780_0007_8007_8000_0F00_0000_0000;
row55<=512'h0000_7038_0000_FFF0_0E00_003F_FFFF_FFC0_0000_0000_0000_0000_0300_0000_007F_FC00_01F8_0078_01C0_0780_0007_8007_C000_1FC0_0000_0000;
row56<=512'h0000_7070_0000_7FE0_0400_0007_FFFF_FF80_0000_0000_0000_0000_0600_0000_000F_FC00_03F0_0070_0180_0780_0007_8003_FFFF_FF80_0000_0000;
row57<=512'h0000_7060_0000_0000_0000_0000_3FFF_FF80_0000_0000_0000_0000_0600_0000_0003_F800_03E0_0060_0100_0300_0007_8003_FFFF_FF00_0000_0000;
row58<=512'h0000_7080_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0C00_0000_0000_F000_0000_0000_0000_0200_0007_8000_FFFF_FE00_0000_0000;
row59<=512'h0000_7100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1800_0000_0000_E000_0000_0000_0000_0000_0007_8000_0000_0000_0000_0000;
row60<=512'h0000_4000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0007_0000_0000_0000_0000_0000;
row61<=512'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0004_0000_0000_0000_0000_0000;
row62<=512'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
row63<=512'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
end
5'b10000:begin
row0<=512'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
row1<=512'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
row2<=512'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_4000_0800_0000;
row3<=512'h0000_0000_0000_0000_0000_0000_0400_0000_0000_001C_0000_0000_0000_0200_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0002_0000_0000_0000_E000_0E00_0000;
row4<=512'h0000_0000_0000_0000_0000_0000_0E00_0000_0000_001F_0000_0000_0000_0380_0C00_0000_0000_0000_0000_0000_0000_0000_0000_0800_0000_0003_8000_0000_0000_F800_0F00_0000;
row5<=512'h0000_0000_0000_0000_0000_0000_0F80_0000_0000_003F_0000_0000_0000_03F0_0F00_0000_0000_0000_0000_0000_000C_0000_0000_1C00_0000_0003_F000_0000_0000_FC00_1FC0_0000;
row6<=512'h0000_0000_0000_0000_0000_0000_0F80_0000_0000_003E_0000_0000_0000_03E0_0FC0_0000_0000_0000_0000_0000_000F_FFFF_FFFF_FF00_0000_0003_E000_0000_0001_F000_1F80_0000;
row7<=512'h0000_0000_0000_0000_0000_0100_0F00_0000_0000_003C_0000_0000_0000_03C0_0F00_0000_0000_0000_0000_0000_000F_FFFF_FFFF_FF00_0000_0003_C000_0000_0001_F000_1F00_0000;
row8<=512'h0000_0000_0000_0000_0180_0180_1E00_0000_0000_0038_0000_0000_0000_0380_0F00_0000_0000_0000_0000_0000_000E_0000_0000_1E00_0000_0003_C000_0000_0001_E000_3F80_0000;
row9<=512'h0000_0000_0000_0000_01FF_FFE0_1E00_0800_0000_0070_0000_0000_0000_0380_0F00_0000_0000_0000_0000_0000_000E_0000_0000_1C00_0000_0003_C000_0000_0001_E000_3C80_0000;
row10<=512'h0000_0000_0000_0000_01FF_FFE0_1C00_1C00_0000_0070_0000_0000_0000_0380_0F00_0000_0000_0000_0000_0000_000E_0001_C000_1C00_0000_0003_C000_0000_0003_C000_7CC0_0000;
row11<=512'h0000_0000_0000_0000_01E0_0380_3FFF_FE00_0000_0060_0000_0000_0000_0380_0F00_0000_0000_0000_0000_0000_000E_0001_F000_1C00_0000_0003_C000_0400_0003_C000_7840_0000;
row12<=512'h0000_0000_0000_0000_01E0_0380_3FFF_FF00_0040_00E0_0000_0400_0000_0380_0F00_0000_0000_0000_0000_0000_000E_0001_E000_1C00_0000_0003_C000_0E00_0003_8000_7860_0000;
row13<=512'h0000_0000_0000_0000_01E0_0380_3800_3E00_0060_00C0_0000_0E00_0000_0380_0F00_0000_0000_0000_0000_0000_000E_0001_C000_1C00_0000_0003_C000_1F00_0007_8000_F030_0000;
row14<=512'h0000_0000_0000_0000_01E0_0380_7800_3C00_007F_FFFF_FFFF_FF80_0000_0380_0F00_0000_0000_0000_0000_0000_000E_0001_C000_1C00_07FF_FFFF_FFFF_FF80_0007_0000_F030_0000;
row15<=512'h0000_0000_0000_0000_01E0_0380_7000_7800_007F_FFFF_FFFF_FF80_0000_0380_0F00_0000_0000_0000_0000_0000_000E_0001_C000_1C00_03FF_FFFF_FFFF_FFC0_000F_0001_E018_0000;
row16<=512'h0000_0000_0000_0000_01E0_0380_6800_7800_0078_0000_0000_0F00_0000_0380_0F00_0000_0000_0000_0000_0000_000E_0001_C060_1C00_0100_001F_D000_0000_000F_0001_E01C_0000;
row17<=512'h0000_0000_0000_0000_01E0_0380_EC00_F000_0078_0000_0000_0E00_0000_0380_0F00_0300_0000_0000_0000_0000_000E_0001_C0F0_1C00_0000_001F_D800_0000_000E_0003_C00E_0000;
row18<=512'h0000_0000_0000_0000_01E0_0380_CC01_E000_0078_0000_0000_0E00_0000_0380_0F00_0780_0000_0000_0000_0000_000E_0FFF_FFF8_1C00_0000_003F_CC00_0000_001E_0003_800F_0000;
row19<=512'h0000_0000_0000_0000_01E0_0381_C601_E000_0078_0000_0000_0E00_0000_0380_0F00_0FC0_0000_0000_0000_0000_000E_07FF_FFFC_1C00_0000_007F_CC00_0000_001C_0007_8007_8000;
row20<=512'h0000_0000_0000_0000_01E0_0381_8703_C000_0078_0000_0000_0E00_0000_0380_0F00_1FE0_0000_0000_0000_0000_000E_0201_C000_1C00_0000_007B_C600_0000_003F_000F_0003_C000;
row21<=512'h0000_0000_0000_0000_01E0_0383_8303_C000_0078_0000_0000_0E00_0FFF_FF80_0F00_3F80_0000_0000_0000_0000_000E_0001_C000_1C00_0000_00F3_C700_0000_003F_C00E_0003_E000;
row22<=512'h0000_0000_0000_0000_01E0_0383_0387_8000_0078_0000_0000_0E00_07FF_FF80_0F00_FC00_0000_0000_0000_0000_000E_0001_C000_1C00_0000_01E3_C380_0000_0077_C01E_0001_F000;
row23<=512'h0000_0000_0000_0000_01FF_FF86_01CF_0000_0078_0000_0000_0E00_0000_0380_0F01_F000_0000_0000_0000_0000_000E_0001_C000_1C00_0000_03E3_C1C0_0000_0077_801C_0000_FC00;
row24<=512'h0000_0000_0000_0200_01FF_FF86_00EE_0000_0078_0000_0080_0E00_0000_0380_0F03_C000_0000_0000_0000_0000_000E_0001_C000_1C00_0000_03C3_C1C0_0000_00E7_8038_0000_7E00;
row25<=512'h0000_0000_0000_0700_01E1_C38C_00FE_0000_0078_0600_01C0_0E00_0000_0380_0F0F_0000_0000_0000_0000_0000_000E_0001_C00C_1C00_0000_0783_C0F0_0000_00C7_8070_0000_3F80;
row26<=512'h0000_0000_0000_0F80_01E1_C308_007C_0000_0078_07FF_FFE0_0E00_0000_0380_0F1C_0000_0000_0000_0000_0000_000E_0001_C01E_1C00_0000_0F03_C078_0000_01C7_80E0_0000_1FF0;
row27<=512'h0000_0000_0000_1FC0_0181_C010_007C_0000_0078_07FF_FFF0_0E00_0000_0380_0F70_0000_0000_0000_0000_0000_000E_FFFF_FFFF_1C00_0000_1E03_C03C_0000_0187_80C4_0000_0FF8;
row28<=512'h1FFF_FFFF_FFFF_FFE0_0001_C000_00FE_0000_0078_0780_01E0_0E00_0000_0380_0FC0_0000_0000_0000_0000_0000_000E_7FFF_FFFF_9C00_0000_3C03_C03F_0000_0307_8187_0000_07C0;
row29<=512'h0FFF_FFFF_FFFF_FFF0_0001_C000_01FF_8000_0078_0780_01C0_0E00_0000_0380_0F00_0000_0000_0000_0000_0000_000E_3000_0000_1C00_0000_7803_C01F_8000_0707_8307_C000_0300;
row30<=512'h0600_0000_0000_0000_0001_C000_03EF_C000_0078_0780_01C0_0E00_0000_0380_0F00_0000_0000_0000_0000_0000_000E_0000_0000_1C00_0000_F003_C00F_F000_0607_8607_C001_0000;
row31<=512'h0000_0000_0000_0000_0001_C000_07C3_F000_0078_0780_01C0_0E00_0000_0380_0F00_0000_0000_0000_0000_0000_000E_0000_0000_1C00_0001_E003_C003_FC00_0C07_8C07_8003_8000;
row32<=512'h0000_0000_0000_0000_0101_C100_0F81_FC00_0078_0780_01C0_0E00_0000_0380_0F00_0000_0000_0000_0000_0000_000E_0000_0000_1C00_0003_8003_C001_FFC0_1807_9807_8007_C000;
row33<=512'h0000_0000_0000_0000_01C1_C380_1E00_FF00_0078_0780_01C0_0E00_0000_0380_0F00_0000_0000_0000_0000_0000_000E_0200_0040_1C00_000F_0003_C000_FFF8_1007_A007_800F_E000;
row34<=512'h0000_0000_0000_0000_01F1_FFC0_3C00_7FE0_0078_0780_01C0_0E00_0000_0380_0F00_0000_0000_0000_0000_0000_000E_0180_00E0_1C00_001C_0003_C000_3FC0_0007_8007_801F_F000;
row35<=512'h0000_0000_0000_0000_01E1_FFE0_7800_1FFC_0078_0780_01C0_0E00_0000_0380_0F00_0000_0000_0000_0000_0000_000E_01FF_FFF0_1C00_0038_0003_C000_0F80_0007_8007_803F_0000;
row36<=512'h0000_0000_0000_0000_01C1_C000_F000_1FF0_0078_0780_01C0_0E00_0000_0380_0F00_0000_0000_0000_0000_0000_000E_01FF_FFF8_1C00_00E0_0003_C000_0300_0007_8007_807C_0000;
row37<=512'h0000_0000_0000_0000_01C1_C003_F000_3BC0_0078_0780_01C0_0E00_0000_0380_0F00_0000_0000_0000_0000_0000_001E_01C0_00E0_1C00_01C0_0003_C000_0000_0007_8007_81F0_0000;
row38<=512'h0000_0000_0000_0000_01C1_C007_FFFF_FC80_0078_0780_01C0_0E00_0000_0380_0F00_0000_0000_0000_0000_0000_001E_01C0_00E0_1C00_0700_0003_C000_0000_0007_8007_83C0_0000;
row39<=512'h0000_0000_0000_0000_01C1_C01E_7FFF_FE00_0078_0780_01C0_0E00_0000_0380_0F00_0000_0000_0000_0000_0000_001C_01C0_00E0_1C00_1C00_0003_8000_0000_0007_8007_8F00_0000;
row40<=512'h0000_0000_0000_0000_01C1_C038_7800_3C00_0078_0780_01C0_0E00_0000_0380_0F00_0000_0000_0000_0000_0000_001C_01C0_00E0_1C00_0000_0002_0000_0000_0007_8007_9C00_0000;
row41<=512'h0000_0000_0000_0000_01C1_C0E0_7800_3800_0078_07FF_FFC0_0E00_0000_0380_0F00_0080_0000_0000_0000_0000_001C_01C0_00E0_1C00_0000_0000_0000_0000_0007_8007_F000_0000;
row42<=512'h0000_0000_0000_0000_01C1_C100_7800_3800_0078_07FF_FFC0_0E00_0000_0380_0F00_0080_0000_0000_0000_0000_001C_01C0_00E0_1C00_0000_0000_0000_0000_0007_8007_C000_0000;
row43<=512'h0000_0000_0000_0000_01C1_C000_7800_3800_0078_0780_01C0_0E00_0000_0380_0F00_0080_0000_0000_0000_0000_003C_01C0_00E0_1C00_0000_0000_0000_0000_0007_8007_8000_0000;
row44<=512'h0000_0000_0000_0000_01C1_C000_7800_3800_0078_0780_01C0_0E00_0000_0F80_0F00_0080_0000_0000_0000_0000_0038_01C0_00E0_1C00_0004_0000_0001_0000_0007_8007_8000_0600;
row45<=512'h0000_0000_0000_0000_01C1_C000_7800_3800_0078_0780_01C0_0E00_0000_7B80_0F00_0080_0000_0000_0000_0000_0038_01C0_00E0_1C00_0004_0200_1000_C000_0007_8007_8000_0600;
row46<=512'h0000_0000_0000_0000_01C1_C000_7800_3800_0078_0780_0180_0E00_0003_E380_0F00_00C0_0000_0000_0000_0000_0038_01FF_FFE0_1C00_000C_0300_1800_E000_0007_8007_8000_0600;
row47<=512'h0000_0000_0000_0000_01C1_C000_7800_3800_0078_0600_0000_0E00_003F_8380_0F00_00C0_0000_0000_0000_0000_0070_01FF_FFE0_1C00_000C_0380_0E00_7000_0007_8007_8000_0600;
row48<=512'h0000_0000_0000_0000_01C1_C1F0_7800_3800_0078_0000_0000_0E00_03FE_0380_0F00_00C0_0000_0000_0000_0000_0070_01C0_00E0_1C00_000C_01C0_0F00_3800_0007_8007_8000_0600;
row49<=512'h0000_0000_0000_0000_01C1_DF80_7800_3800_0078_0000_0000_0E00_0FF8_0380_0F00_01C0_0000_0000_0000_0000_0060_01C0_00E0_1C00_001C_01E0_0780_3E00_0007_8007_8000_0600;
row50<=512'h0000_0000_0000_0000_01C1_FC00_7800_3800_0078_0000_0000_0E00_0FE0_0380_0F00_01C0_0000_0000_0000_0000_00E0_01C0_00F0_1C00_001C_00E0_07C0_1F00_0007_8007_8000_0600;
row51<=512'h0000_0000_0000_0000_01DF_E000_7800_3800_0078_0000_0000_0E00_0780_0380_0F00_01C0_0000_0000_0000_0000_00C0_01C0_0080_1C00_003C_00F0_03C0_1F00_0007_8007_8000_0600;
row52<=512'h0000_0000_0000_0000_01FF_0000_7800_3800_0078_0000_0000_0E00_0300_0380_0F00_01E0_0000_0000_0000_0000_01C0_0100_0000_1C00_007C_00F8_03E0_0F80_0007_8007_8000_0E00;
row53<=512'h0000_0000_0000_0000_1FFC_0000_7800_3800_0078_0000_0000_1E00_0200_0380_0F00_03F0_0000_0000_0000_0000_0180_0000_0000_1C00_0078_0078_03E0_0F80_0007_8007_8000_0E00;
row54<=512'h0000_0000_0000_0000_0FE0_0000_7FFF_F800_0078_0000_007F_FE00_0000_0380_0F80_07F0_0000_0000_0000_0000_0380_0000_0000_3C00_00F8_0078_03E0_0780_0007_8007_8000_0F00;
row55<=512'h0000_0000_0000_0000_0F80_0000_7FFF_F800_0078_0000_001F_FE00_0000_0380_07FF_FFF0_0000_0000_0000_0000_0300_0000_007F_FC00_01F8_0078_01C0_0780_0007_8007_C000_1FC0;
row56<=512'h0000_0000_0000_0000_0600_0000_7800_3800_0078_0000_0003_FE00_0000_0380_07FF_FFE0_0000_0000_0000_0000_0600_0000_000F_FC00_03F0_0070_0180_0780_0007_8003_FFFF_FF80;
row57<=512'h0000_0000_0000_0000_0000_0000_7800_3800_0078_0000_0000_FC00_0000_0380_01FF_FF00_0000_0000_0000_0000_0600_0000_0003_F800_03E0_0060_0100_0300_0007_8003_FFFF_FF00;
row58<=512'h0000_0000_0000_0000_0000_0000_7800_3800_0078_0000_0000_7800_0000_03C0_0000_0000_0000_0000_0000_0000_0C00_0000_0000_F000_0000_0000_0000_0200_0007_8000_FFFF_FE00;
row59<=512'h0000_0000_0000_0000_0000_0000_7800_3800_0070_0000_0000_7000_0000_0200_0000_0000_0000_0000_0000_0000_1800_0000_0000_E000_0000_0000_0000_0000_0007_8000_0000_0000;
row60<=512'h0000_0000_0000_0000_0000_0000_7000_2000_0040_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0007_0000_0000_0000;
row61<=512'h0000_0000_0000_0000_0000_0000_4000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0004_0000_0000_0000;
row62<=512'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
row63<=512'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
end
endcase
end
end
endmodule
